package id_pkg;
    typedef enum logic[3:0] { 
        STORE = 4'b0111,
        NOP = 4'b1111
    } cpu_instructions;
endpackage : id_pkg