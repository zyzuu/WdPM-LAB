module top()
    
endmodule : top