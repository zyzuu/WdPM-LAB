module alu_accumulator_tb();
    
endmodule : alu_accumulator_tb