module simple_top(
    input clk
);
    
endmodule : simple_top