`ifndef opcodes
`define opcodes

`define ADD 0000;
`define SUBTRACT 0001;
`define AND_OP 0010;
`define OR_OP 0011;
`define XOR_OP 0100;
`define NOT_OP 0101;
`define LOAD 0110;
`define STORE 0111;
`define NOP 1111;
`endif opcodes